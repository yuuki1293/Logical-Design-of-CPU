`timescale 1ps/1ps

// |---|----|------|------|-------|
// | A |  B |  CIN |  Q   |  COUT |
// |---|----|------|------|-------|
// | 0 |  0 |  0   |    0 |  0    |
// |---|----|------|------|-------|
// | 0 |  0 |  1   |    1 |  0    |
// |---|----|------|------|-------|
// | 0 |  1 |  0   |    1 |  0    |
// |---|----|------|------|-------|
// | 0 |  1 |  1   |    0 |  1    |
// |---|----|------|------|-------|
// | 1 |  0 |  0   |    1 |  0    |
// |---|----|------|------|-------|
// | 1 |  0 |  1   |    0 |  1    |
// |---|----|------|------|-------|
// | 1 |  1 |  0   |    0 |  1    |
// |---|----|------|------|-------|
// | 1 |  1 |  1   |    1 |  1    |
// |---|----|------|------|-------|

module fulladd_tp;

reg A, B, CIN;
wire Q, COUT;

// シミュレーションステップの設定
parameter STEP = 100000;

// テスト対象インスタンス
fulladd fulladd(A, B, CIN, Q, COUT);

// テスト入力
initial begin
    // VCDファイル出力
    $dumpfile("fulladd.vcd");
    $dumpvars(0, fulladd_tp);

          A = 1'b0; B = 1'b0; CIN = 1'b0; // 0 + 0 + 0 -> Q = 0, COUT = 0
    #STEP A = 1'b0; B = 1'b0; CIN = 1'b1; // 0 + 0 + 1 -> Q = 1, COUT = 0
    #STEP A = 1'b0; B = 1'b1; CIN = 1'b0; // 0 + 1 + 0 -> Q = 1, COUT = 0
    #STEP A = 1'b0; B = 1'b1; CIN = 1'b1; // 0 + 1 + 1 -> Q = 0, COUT = 1
    #STEP A = 1'b1; B = 1'b0; CIN = 1'b0; // 1 + 0 + 0 -> Q = 1, COUT = 0
    #STEP A = 1'b1; B = 1'b0; CIN = 1'b1; // 1 + 0 + 1 -> Q = 0, COUT = 1
    #STEP A = 1'b1; B = 1'b1; CIN = 1'b0; // 1 + 1 + 0 -> Q = 0, COUT = 1
    #STEP A = 1'b1; B = 1'b1; CIN = 1'b1; // 1 + 1 + 1 -> Q = 1, COUT = 1
    #STEP $finish;
end

// コンソール出力
initial $monitor($stime, " A=%b B=%b CIN=%b Q=%b COUT=%b", A, B, CIN, Q, COUT);

endmodule